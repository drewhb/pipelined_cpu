module hazardunit(IFIDWrite,PCWrite,HazardMux);

   output     IFIDWrite, PCWrite, HazardMux;
   
   
   assign IFIDWrite = 1;
   assign PCWrite = 1;
   assign HazardMux = 0;
   
endmodule
